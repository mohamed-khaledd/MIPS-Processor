module DataMemory(
    input clk,
    input [31:0] addr,
    input [31:0] write_data,
    input write_enable,
    output [31:0] read_data
);

  /* Module Description:
     - The module has 4 inputs:
       1) addr, which is the address of the data to be read.
       2) write_data, which is the data to be written in the data memory.
       3) clk, which is the clock signal.
       4) write_enable, which is the write enable signal.
     - The module has an output read_data which is the data read.
  */
  
    reg [31:0] memory [0:4095];
    integer i;

    initial begin
        for (i = 0; i < 4096; i = i + 1) begin
            memory[i] = 32'b0;    // // Initializing all memory to zero
        end
    end

    assign read_data = memory[addr[31:2]];

    always @(posedge clk) begin
        if (write_enable)
            memory[addr[31:2]] <= write_data;
    end
endmodule
